module game(input clk, input rst, input [3:0]choice, output reg [1343:0] frame);

reg[4:0]S;
reg[4:0]NS;
reg[4:0]LS;
reg[7:0]selection;

always@(posedge clk or negedge rst)
begin
    if (rst == 1'b0)
    begin
        S <= START;
    end
    else
        S <= NS;
end

reg userInput;

parameter START = 5'd0,
          START_2 = 5'd1,
          EXAM = 5'd2,
          NOW = 5'd3,
          NOW_2 = 5'd4,
          PRINT = 5'd5,
			 FOOD = 5'd6,
			 SINK = 5'd7,
			 FIRE = 5'd8,
			 PUT_OUT = 5'd9,
			 GIVE_UP = 5'd10,
			 ALT_NOW = 5'd11,
			 NO_PRINT = 5'd12,
			 ALIVE = 5'd13,
			 DEAD = 5'd14,
			 NO_FOOD = 5'd15,
			 TWO_DAYS = 5'd16,
			 ONE_DAY = 5'd17,
			 ZERO_DAYS = 5'd18,
			 PRESSURE = 5'd19,
			 SURPRISE = 5'd20,
			 CRUMBLE = 5'd21,
			 GAMER = 5'd22,
			 NEVER = 5'd23,
          confirmInput = 5'd24;

always@(*)
begin
    case(S)
        START: 
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = START;
        end
        START_2:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = START_2;
        end
        EXAM:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = EXAM;
        end
        NOW:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = NOW;
        end
        NOW_2:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = NOW_2;
        end
        PRINT:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = PRINT;
        end
		  FOOD:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = FOOD;
        end
		  SINK:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = SINK;
        end
		  FIRE:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = FIRE;
        end
		  PUT_OUT:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = PUT_OUT;
        end
		  GIVE_UP:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = GIVE_UP;
        end
		  ALT_NOW:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = ALT_NOW;
        end
		  NO_PRINT:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = NO_PRINT;
        end
		  ALIVE:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = ALIVE;
        end
		  DEAD:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = DEAD;
        end
		  NO_FOOD:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = NO_FOOD;
        end
		  TWO_DAYS:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = TWO_DAYS;
        end
		  ONE_DAY:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = ONE_DAY;
        end
		  ZERO_DAYS:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = ZERO_DAYS;
        end
		  PRESSURE:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = PRESSURE;
        end
		  SURPRISE:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = SURPRISE;
        end
		  CRUMBLE:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = CRUMBLE;
        end
		  GAMER:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = GAMER;
        end
		  NEVER:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = NEVER;
        end
        confirmInput:
        begin
            if (userInput == 1'b0)
            begin
                case(LS)
                    START:
						  begin
						      NS = START_2;
						  end
                    START_2:
						  begin
						      NS = EXAM;
						  end
						  EXAM:
						  begin
								case(selection)
                                    8'd1: NS = NOW;
                                    8'd2: NS = TWO_DAYS;
                                    8'd3: NS = NEVER;
                                    8'd4: NS = EXAM;
                                    default: NS = confirmInput;
                                endcase
						  end
						  NOW:
						  begin
						      NS = NOW_2;
						  end
						  NOW_2:
						  begin
                                case(selection)
                                    8'd1: NS = NO_PRINT;
                                    8'd2: NS = PRINT;
                                    8'd3: NS = NO_PRINT;
                                    8'd4: NS = PRINT;
                                    default: NS = confirmInput;
                                endcase
						  end
						  PRINT:
						  begin
                                case(selection)
                                    8'd1: NS = FOOD;
                                    8'd2: NS = NO_FOOD;
                                    8'd3: NS = FOOD;
                                    8'd4: NS = NO_FOOD;
                                    default: NS = confirmInput;
                                endcase
						  end
						  FOOD:
						  begin
                                case(selection)
                                    8'd1: NS = SINK;
                                    8'd2: NS = PUT_OUT;
                                    8'd3: NS = SINK;
                                    8'd4: NS = PUT_OUT;
                                    default: NS = confirmInput;
                                endcase
						  end
						  SINK:
						  begin
						      NS = FIRE;
						  end
						  FIRE:
						  begin
						      NS = FIRE;
						  end
						  PUT_OUT:
						  begin
                                case(selection)
                                    8'd1: NS = ALT_NOW;
                                    8'd2: NS = GIVE_UP;
                                    8'd3: NS = PUT_OUT;
                                    8'd4: NS = PUT_OUT;
                                    default: NS = confirmInput;
                                endcase
						  end
						  GIVE_UP:
						  begin
						      NS = GIVE_UP;
						  end
						  ALT_NOW:
						  begin
                                case(selection)
                                    8'd1: NS = PRINT;
                                    8'd2: NS = NO_PRINT;
                                    8'd3: NS = PRINT;
                                    8'd4: NS = NO_PRINT;
                                    default: NS = confirmInput;
                                endcase
						  end
						  NO_PRINT:
						  begin
                                case(selection)
                                    8'd1: NS = DEAD;
                                    8'd2: NS = ALIVE;
                                    8'd3: NS = DEAD;
                                    8'd4: NS = ALIVE;
                                    default: NS = confirmInput;
                                endcase
						  end
						  ALIVE:
						  begin
						      NS = ALIVE;
						  end
						  DEAD:
						  begin
						      NS = DEAD;
						  end
						  NO_FOOD:
						  begin
						      NS = NO_FOOD;
						  end
						  TWO_DAYS:
						  begin
                                case(selection)
                                    8'd1: NS = ONE_DAY;
                                    8'd2: NS = NOW;
                                    8'd3: NS = TWO_DAYS;
                                    8'd4: NS = TWO_DAYS;
                                    default: NS = confirmInput;
                                endcase
						  end
						  ONE_DAY:
						  begin
                                case(selection)
                                    8'd1: NS = ZERO_DAYS;
                                    8'd2: NS = NOW;
                                    8'd3: NS = ONE_DAY;
                                    8'd4: NS = ONE_DAY;
                                    default: NS = confirmInput;
                                endcase
						  end
						  ZERO_DAYS:
						  begin
                                case(selection)
                                    8'd1: NS = GAMER;
                                    8'd2: NS = PRESSURE;
                                    8'd3: NS = ZERO_DAYS;
                                    8'd4: NS = ZERO_DAYS;
                                    default: NS = confirmInput;
                                endcase
						  end
						  PRESSURE:
						  begin
                                case(selection)
                                    8'd1: NS = CRUMBLE;
                                    8'd2: NS = SURPRISE;
                                    8'd3: NS = PRESSURE;
                                    8'd4: NS = PRESSURE;
                                    default: NS = confirmInput;
                                endcase
						  end
						  SURPRISE:
						  begin
						      NS = SURPRISE;
						  end
						  CRUMBLE:
						  begin
						      NS = CRUMBLE;
						  end
						  GAMER:
						  begin
						      NS = GAMER;
						  end
						  NEVER:
						  begin
						      NS = NEVER;
						  end
                endcase
            end
            else
                NS = confirmInput;
        end
    endcase
end

always@(posedge clk or negedge rst)
begin
    if (rst == 1'b0)
	 begin
        frame <= 1344'b011000000001000001011000001000011100001100000010001111111000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110000000011100001000001101100011000110000001110001010010001100010010000010000001001000110100010110001101000110000111100100010000100001001000100101000110000000000011010011000100011000000010010100001001100100110001110000110100100110001110100011000000100001110000110100100110001000000110100101000000100011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000101;
        LS <= START;
	 end
    else
	 begin
        case(S)
            START:
            begin
                frame <= 1344'b011000000001000001011000001000011100001100000010001111111000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110000000011100001000001101100011000110000001110001010010001100010010000010000001001000110100010110001101000110000111100100010000100001001000100101000110000000000011010011000100011000000010010100001001100100110001110000110100100110001110100011000000100001110000110100100110001000000110100101000000100011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000101;
                LS <= START;
            end
            START_2:
            begin
                frame <= 1344'b010111000100100000100100011000100110000111000010010001100000001001010000100110010011000111000011010010010100011000011100001101100011000100110000111000010010001100000001000111000000000010001000001110001100010011000111010001100001100000000000010100000100100011000110000001110001010000100011000110100011010001101000110100011010001101000110001001000001000001011000010000000100010011000100000011100001101011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100101101000011100001001000110000111000100010000011000010000100011000110000111000001011000110001001100001110000100000000100101000010011001001100011100001101001001010001100001000001001010001100000000001001010001101000110100011000001010001110000101100010110001110001011000100101000110000010100100010001110000110010001101000110100011010001100001011000010000001010010011100011000100110001110100011000100010001000000011000001110010011100011010001101000110011100010001100110111100011001101101000110011010110001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000101;
                LS <= START_2;
            end
				EXAM:
            begin
                frame <= 1344'b011001000011100010100100011000000000010001000010010001100001111000101100000000011000000100000011010000110100011000000100001110001010000011010010011000010000100010010010001001100100010001000000101000001001000110011011010001100010110000011100001000001101100011000110000001110001010010001100010001000010000000100000100000100000101010000100000000000011011000110001111000011000000000000100000010111000110000010100100010001110000110010001101000110100011000111010010001011111010001100100011000000000011000001000000010000100100001110000110101111101000110010001000100110001000001001010001100010011000011100001001000110011011001111000111011100011000001000010111000000000011000111111100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110011010110001100011101000111010001100001000001001110001100001101000111000101101000110100011010001101000110100011001101101000110001110100011101000110000100000100111000110000101100000000010011000010000100011000110100011010001100110111100011000111010001110100011000010000010011100011000011010000100001010100001000010001100011010001101000110;
                LS <= EXAM;
            end
				NOW:
            begin
                frame <= 1344'b011001000011100010100100011000000110000100000001000010000000011000010010001100010011000111010001100000001000010000100010000100001001000011110001110000110100100100001000000000100010110000100100011000000000001101000001110001100010010001001100000000010001001001110001100010011000011100001001000110000010000101110000000000110001111101000110001101000100101000110001100000011100010100100011000010110001110000000000000111000110001001100001110000100100011000001010001000000101100001001000010100011000110000001110001010010001100010010000010000001001000110100011010001100011000000111000101000010001100011000011110010001000100000011010010011000010000100010111110100011001000100010011000011100000000010010100011000000010000100000010000011011000110000000010001100010110000011100010000001011000010000100100001000000110100000100000100100011000010000010011100000100100101000110000101100000000010010001001110001100010100001001000001000111110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000101;
                LS <= NOW;
            end
				NOW_2:
            begin
                frame <= 1344'b001110100011101000110001100000011100010100100011000011110010001000100000011010010011100011000011100010100001001100100110000111000010010001100000100001011100000000001100100000010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110011010110001100100111000111010000101000110010001010000010001100100011000011010001110001001110001100000000100011010001101000110000001000000000010101000010000011000000000000110101111111000110100011010001101000110100011010001100110110100011001100100000100001001010000101000110001001100001110000100100011010001101000110100011010001101000110100011010001100001111001000100010000001101001001100001000010001100011000011000010100001001000100111000110100011010001101000110000000100001001000110001010000100100000100000001101111101000110100011010001101000110100011010001100110111100011001001110001110100001010001100001000000110100010101000110000100000100101000110001001100011100001110100011010001100000100001011100011110000100000110100100100001000001010100001000111111100011010001101000110100011001110001000110011001000001000010010100001010001100001010000100000010110001011100011000100100001110000110000001001000110100011000100110010001000010000001000010010011111110001101000110100011010001101000110100011010001101000110;
                LS <= NOW_2;
            end
				PRINT:
            begin
                frame <= 1344'b011001000011100010100100011000011110010001000100000011010010011100011000011100010100001001110001101000110100011000100110000111000010010001100000100001011100000000001100100001010001100000001001010000100111000110100011010001100000000001000100001001000110001001000011100001110000110110001101000110100011010001101000110100011010001101000110001000100001000001100000100000011010000011000010000000111000110000111000001011000110001100000011100010100001000100001110010100000110100001100000100001000101111101000110001110100011101000110001100000011100010100100011010001100001100000000000010100000100100011000001010001110000111000000111000000100011010001101000110100011010001101000110011010110001100110010000010000100101000010100011000101100001000001001100001111000110100011010001101000110100011010001101000110000001000001110000100000010000100100000100011111010001101000110100011010001101000110100011010001100110110100011001001110001110100001010001100010010000101000010000001111100011000001010001110000111000000111000110011011110001100110010000010000100101000010100011000101100001000001001100001110001110001010000100111000110100011010001101000110000001000001110000100000010000100100000100100011010001101000110100011010001101000110100011010001100111000100011001001110001110100011000100110001000000110000001000111111100011010001101000110100011010001101000110;
                LS <= PRINT;
            end
				FOOD:
            begin
                frame <= 1344'b011001000011100010100100011000001100001110100011000100110001110100011000011000000000000101000001001000110100011000001010001110000111000000111000010100011000000010010100001001110001101000110100011010001101000110100011010001100000000000001000000100001000000001100001000001101001001100000000001011000101100110001000110001001000001000010011001001100001110000100100011000001000010111000000000011001000110000111000011011000110100011010001101000110100011000001010001000001000100001000111111100011001100000000111000000000100111000110000001100011101000110100011010001100011000000111000101001000110000001100011101000000100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011001101011000110010100100000000001101000100000000100111111100011010001101000110100011010001101000110100011010001100110110100011001011000010011000000000110001000110000001000000000001011000110001111111000110100011010001101000110011011110001100101101000011100100010001110001011010001100010011000011100001001000110000010000101110000000000110010001101000110000100000011011000110001001100001110000100100011000100100001000000110100010100111111100011010001100111000100011001010010010100001001110001100001000001001110001100001110001010000100110111111100011010001101000110;
                LS <= FOOD;
            end
				SINK:
            begin
                frame <= 1344'b011001000011100010100100011000100110000111001000100011100010110100011000100110000111000010010001101000110100011000001000010111000000000011001000110000100000011011000110001001100001110000100100011000100100001000000110100010100010011000011100010000001101000101000010000001101000011010001100001000001001110001100010110000100000010110001011000101100000000001101000001110001100001000000110110001100010110000000000100110000100001000101111101000110100011001100100001110001010010001100000000001000100001001000110001011000100010001110000110100001100111110100011010001100100010001001110001100001011000000000011010000011001001010001100001000000110110001100000000100011010001101000110000111100011100010011100011000011100000101100011000001110001110001001110001100001110000100000010111000110100011000010000001101001001000100110000100000000000000110111110100011001100100001110001010000100011000110100011010001100001010000100000100110000010000011100001000001101100011000001100001110000010000100101000110001010000011111000110000100000011011000110000010100010110000000000110000001000010010100011000000000001101000001110001101000110100011000100110000111000010010001100000101000100000100010000100100011000100000010100000100000000100001010000101100110000010010000111100100010000100000000000000110010010011111010001101000110100011010001101000110100011010001101000101;
                LS <= SINK;
            end
				FIRE:
            begin
                frame <= 1344'b010110100001110000100100011000001010001000001000100001001000110001001100100010000000001010100001000001011001001000000000000010001000100011100010010001001010001100010011000011100001001000110001010100001000010001001100010001100000101000101100000000001100000110000000000000001000101100001001000110000011000100010000000001001000100100111110010110100001110000100100011000101000001101000100000101010000100001000100100100001000001001100110001000110100011000001110000000001001010001100001101000111010001100000010000011100000000001101000001000001000111110100011010001100110010000111000101001000110000100000011000001100000010000000110001000000000000100110000100000101100110001000110000011000100010000000000001100101000000000001001100001001000110001011000010000010011000011110001100000000100011000000110000100000011000100010000100000010010001100001000000110110001101000110100011010001101000110100011010001100000100000110100001100001000000110100001000000100001000100010000001101000011001111101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000111100000000010010001001000001000000011011111110001100011010100010010001101000110;
                LS <= FIRE;
            end
				PUT_OUT:
            begin
                frame <= 1344'b011001000011100010100100011000001100010001000000000000011000110001001100001110000100100011010001101000110100011000001000010111001001100010000001101000011000101000001000001001000001110000100001000110001100000000000110100000110001111001010000100111000110000111000101000010011100011000100110000111000010010001101000110100011010001101000110000010100010000010001000010001111101000110011001000011100010100100011000011010000100000010000000111000110000000000011010000100001011010001100000100001011100000000001100100001010001100000001001010000100111000110100011010001100000010000000000011011000001001001110001100000111000010000010110001111100011000000010010100001001110001101000110001000000101000000100001001000100110001000000111000011011000110000100000001011000110000100000100111000001001001000101100001110001000100100110000111100011000010000010011011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011001101011000110010000000001000010011100011000011010000100001011010001100000100001011100000000001100100011010001100110110100011001001110001110001001110001100010110000111000100010010011000011110001100001000001001110001101000110;
                LS <= PUT_OUT;
            end
				GIVE_UP:
            begin
                frame <= 1344'b011001000011100010100100011000100110000111000100000011010001010100011000110000001110001010010001101000110100011000011000000000000001100001001000110000000010001100000110000111000011100000011100011010001101000110100011010001100000100000010100001010001110001000100100111000110000000000001010010011000010000100011000110100011010001101000110000000000010110001100000111000100100010011100011000000010010100001000100011010001000000110100001101000110100011000110000001110001010000100011000110000101000010000010011000001000001110000100000110110001101000110100011010001100000011000111000101100001101011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011000111010010001011111010001100100011000000000011000001000000010000100100001110000110110001101000110100011010001100000011000111000001000010010100011000011010001110001001110001100000000000011000100010000100000010001111101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000010100000000001000000101100001000000011011111010001100011111100011010001101000110;
                LS <= GIVE_UP;
            end
				ALT_NOW:
            begin
                frame <= 1344'b011001000011100010100100011000001100001110100011000100110001110100011000001100000100001001110001100000000100011000011010000100001011010001100000100001011100000000001100011111010001100011010001001010001100011000000111000101000000011000111010000101000110001100000011100010100100011000100100000100000010010001100011000000111000101000010001000111100100010001000000110100100110000100001000101111101000110001110100011101000110001100000011100010100100011000011110010001000100000011010010011100011000000000001101000111000100110000111000010000100011000110100011010001100000010000111000011110011000100000010001101000110100011010001101000110100011010001101000110100011010001101000110011010110001100110010000010000100101000010100011001000101000110000101100001000000000001000100011010000100000001110001101000110000110100011100010011000011100010000001101000011001111111000110100011010001101000110100011010001100110110100011001001110001110100001010001100001101000111000100111000110000000000001100000000000100000011011000110011011110001100110010000010000100101000010100011000100110000111000000000100111000110001011000000000010010100011010001101000110000010100101000001101011111110001101000110100011010001101000110100011010001101000110100011010001100111000100011001001110001110100001010001100000110000111010001100000011000100000001100001000001001100000000001011;
                LS <= ALT_NOW;
            end
				NO_PRINT:
            begin
                frame <= 1344'b011001000011100010100100011000001100001110100011000000110001000000011000010000010011000000000010111000110100011000101100001000001001100001111000110001100000011100010100001000110001100000100001011100000000001100011111010001100110010000111000101001000110000011000001000010011100011000110000001110001010000100011000110100011010001101000110000100001010010000000000001110000101000110000000100101000010011100011000000110001000000001110001101000110100011000110000001110001010010001100000010000011100000000010001000011000001001000110000100000100111000000100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110011010110001100101000000010110001100000010000111000101000010001001001000001000111111100011010001101000110100011001101101000110010011100011101000010100011001000101000110000000000010110010110000000000110000010010100011010001101000110100011000001010001110001000100001100000100001001110001101000110100011010001101000110100011010001101000110011011110001100100111000111010000101000110000100000100111000001001001010001100000011000010000000000000011100011001110001000110010001000100111000110001001000001110001110001010000010110000011100011000000010000100100011010001101000110100011000000100000111000000000100010000110000010000000111000110100011010001101000110100011010001101000110;
                LS <= NO_PRINT;
            end
				ALIVE:
            begin
                frame <= 1344'b011001000011100010100001000110001100001000010100100000000000011100011000010000010010100011010001101000110100011000000000001011000100000101010000100011111010001100110010000111000101001000110000010100010110011000100011010001100010011000011100100010001110001010000001100000111100011000100110000111000010010001100000100001011100000000001100001001100001110001000000110100010100001000000110100001101000110000011100011100010110100011010001101000110100011000001000000000001001000110001000110000100000100111000110000100000100100111110100011010001101000110100011010001100110000000011100010000001011000010010001100011000000111000101001000110000000000100010000100100011010001101000110001000100010000000110000011100100111000010100011000011000001110001000100001001000110001001100010000001100000010000101100001110001010000010110000011100011000001110000000001010100001001000110000000100001000000100000110110001100000001000010000100110010011000010000100010111110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000111100000000010010001001000001000000011011111110001100011010100001110001101000110;
                LS <= ALIVE;
            end
				DEAD:
            begin
                frame <= 1344'b011001000011100010100001000110001100001000010100100000000000011100011000010000010010100011010001101000110100011000000110000100000000000000110111110100011001100100001110001010010001100010110000000000010000010011100011010001100000101000111000100011000110000100000100111000110001001100011101000110000001000001110000000001000100001100000100000000000011010000011100011000100110000111000010000011011000110001001000100110000000001000100100110111110100011001011010000111000010010001100000100001011100100110010001000000010001100010011000100000011000000100100011010001100000001000010000011010000100000010100010000010011001001100001000000011100011000110000001110001010001111101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000111100000000010010001001000001000000011011111110001100011010100011010001101000110;
                LS <= DEAD;
            end
				NO_FOOD:
            begin
                frame <= 1344'b011001000011100010100100011000010000000110000110100011100010001000010010001100011000000111000101000010001100011000001110010100000110100001100000100001000110001100000000000110100000111000110001001100000000001010000010010001100010011000011100001001000110000010000101110000000000110010001100001110000110110001100000000000110110001101000110000010000011000001111001001100110001000110001001000100110001110000110000000000000010000011101111101000110100011000110100010010100011001011000001101000100000000100001010000010000100010010010100011010001101000110100011010001100010110000111000101000001011000001110001100001111001010000100111000110000100000100111000010100011010001101000110001100000011100010100100011000001100000100001001110001100000000100011000010110001000001001100100110001011000010000100100010011001010000011110001000000001110001100010110000011100001000001101100011010001101000110100011010001100011000000111000101001000001001000100001001000110000011100101000001101000011000100010011000011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011001100100001110001010010001100000001000000000100010000100000101100110001000110000111100000000010010001001001111110011101100001110001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110;
                LS <= NO_FOOD;
            end
				TWO_DAYS:
            begin
                frame <= 1344'b011001000011100010100100011000010000000110000110100011100010001000010010001100010011000011100001001000110100011000001000010111000000000011001000110000010100011100010001100011000000001000110000001100000000011000011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110010110100001110000100001000100001001000110000000000100010000100100011000011010001110001011010001100110110100011000000110000000001100000100101000110001000100001000001100000000000010000001101000100000011010000110011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110011000000001110000000001001110001100000011000111010001100011000000111000101001000110000001100011101000000100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011001101011000110001110100011101000110000100000100111000110000101100000000010011000010000100011000110100011010001100110110100011000111010001110100011000010000010011100011000011010001110001011010001101000110100011010001101000110;
                LS <= TWO_DAYS;
            end
				ONE_DAY:
            begin
                frame <= 1344'b011001000011100010100100011000010000000110000110100011100010001000010010001100010011000011100001001000110100011000001000010111000000000011001000110000010100011100010001100011000000001000110000001100000000011000011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110010110100001110000100001000100001001000110000100000100101000110000110100011100010110100011001101011000110100011000000110000000001100010001100010001000010000011000000000000100000011010001000000110100001100111110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110011000000001110000000001001110001100000011000111010001100011000000111000101001000110000001100011101000000100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011001101011000110001110100011101000110000100000100111000110000101100000000010011000010000100011000110100011010001100110110100011000111010001110100011000010000010011100011000011010001110001011010001101000110100011010001101000110;
                LS <= ONE_DAY;
            end
				ZERO_DAYS:
            begin
                frame <= 1344'b011001000011100010100100011000010000000110000110100011100010001000010010001100010011000011100001001000110100011000001000010111000000000011001000110000010100011100010001100011000000001000110000001100000000011000011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110010110100001110000100001000100001001000110000000000100010000100100011000011010001110001011010001100110100100011000000110000000001100000100101000110001000100001000001100000000000010000001101000100000011010000110011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110011000000001110000000001001110001100000011000111010001100011000000111000101001000110000001100011101000000100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011001101011000110001110100011101000110000100000100111000110000101100000000010011000010000100011000110100011010001100110110100011000111010001110100011000010000010011100011000011010001110001011010001101000110100011010001101000110;
                LS <= ZERO_DAYS;
            end
				PRESSURE:
            begin
                frame <= 1344'b011001000011100010100100011000001100001110100011000100110001110100011000100100010011000000000100010010011100011000100110000111000010010001100000100001011100000000001100100001010001100000001001010000100111000110100011010001100000010000000000011011000001001001110001100010001000010000011000000100000110000000010000100001000110001101000110000100000001011000110001100000011100010100100011000101100001110001000100010101000110001011000001000001011000101100101000001101000001100001000010001100011000011110010001000010000100100010010001010000100010000100011111010001100011101000111010001100011000000111000101001000000100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110011010110001100100001000111000010110000011100011000011000011000100011000000010000100000010000100011000110100011001101101000110010100000011010000100100011000101100000000001100010001100010011000111010001101000110100011010001101000110100011000001010001000000110100000111000110000111000101000010011100011010001101000110100011010001101000110;
                LS <= PRESSURE;
            end
				SURPRISE:
            begin
                frame <= 1344'b011001000011100010100100011000000110001110100011000101100001110001000100010101000110001011000001000001011000101100101000001101000001100001000010001100011000011110010001000010000100100010010001010000100010000100011111110001100110010000111000101001000110000011000001000010011100011000100110000111000010010001101000110100011010001101000110001011000001110001110000101100001001000110001001100001110001000000110100001101000110000001100011100001101000010000101100001000001001100001111000110011011010001100001100000100000011010010100001001100001000010010100011010001100010011000111010001100010010000111100000000010001000010001111111000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000111100000000010010001001000001000000011011111110001100011011100010010001101000110;
                LS <= SURPRISE;
            end
				CRUMBLE:
            begin
                frame <= 1344'b001110100001000010010000111100010000010011000010010001100010110000011100000000010011100011000110000001110001010000100110000111000100000011010001010100001010001100011000000111000101001000110100011010001101000110100011010001100000010001000100101000001100000000100010110000100100011000101000001101000001100001000010001100011010001101000110000111100100010000100001001000100100010100001000100001000111110100011001000100010011100011010001101000110100011000000100001110001010000010110000011100011000001110000000001010100001001000110000000100001000000100000110110001100010110000111000100010010010000010010001100010011000011100011100010100000011000001110111110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011001001100000000001100000000010000100100011000100100010011000000000100010010011100011010001101000110100011010001100010010000111000011100001101000010000100011000110000110100001000010111001001110001101000110100011010001101000110001001100010000001100000010001111101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000111100000000010010001001000001000000011011111110001100011101100010010001101000110;
                LS <= CRUMBLE;
            end
				GAMER:
            begin
                frame <= 1344'b011001000011100010100100011000011010000100001010100001000010001100011000100110001110000111000010101000110100011000100110000111000010010001100000100001011100000000001100100001010001100000001001010000100111000110100011010001100000001000010000000100000000000110000001001000110000000010001101000110100011010001101000110100011010001101000110000111100100010001110000010100001000010010001001000010000001110000110100000000001011100011000111000101100011011000011110001011000000000110000000100001000110001100010110000100000100110000111100011000000000001011000101110001100010011000011100001001000110000010100100010000100000010010001100010011000100000011000000100100011010001101000110001100000011100010100100011000001110000000000001101111101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000010100000000001000000101100001000000011100011000100110000111000010010001101000110000010000101110000000000110010000101000110000000100101000010011100011000011110000000001001000100100000100000001100000000010011100011000010110001000000010100001000111110100011010001101000110100011010001101000110100011010001100011111100010010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110;
                LS <= GAMER;
            end
				NEVER:
            begin
                frame <= 1344'b011001000011100010100100011000011010000100001010100001000010001100011000100110000000000101000001001000110100011000100110000111000010010001100000100001011100000000001100011111010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001100110010000111000101001000110000010100000000001000000101100001000000011011111010001100011111100011010001101000110;
                LS <= NEVER;
            end
        endcase
    end
end

always@(posedge clk or negedge rst)
begin
    if (rst == 1'b0)
    begin
        userInput <= 1'b0;
        selection <= 1'b0;
    end
    else
    begin
    case(choice)
    4'b1110:
    begin
        userInput <= 1'b1;
        selection <= 8'd1;
    end
    4'b1101:
    begin
        userInput <= 1'b1;
        selection <= 8'd2;
    end
    4'b1011:
    begin
        userInput <= 1'b1;
        selection <= 8'd3;
    end
    4'b0111:
    begin
        userInput <= 1'b1;
        selection <= 8'd4;
    end
    default:
    begin
        userInput <= 1'b0;
        //selection = 8'd0;
    end
    endcase
    end
end

endmodule
