module game(input clk, input rst, input [3:0]choice, output reg [1343:0] frame);

reg[2:0]S;
reg[2:0]NS;
reg[2:0]LS;
reg[7:0]selection;

always@(posedge clk or negedge rst)
begin
    if (rst == 1'b0)
    begin
        S <= START;
    end
    else
        S <= NS;
end

reg userInput;

parameter START = 3'd0,
          firstChoice = 3'd1,
          secondChoice = 3'd2,
          thirdChoice = 3'd3,
          fourthChoice = 3'd4,
          ending       = 3'd5,
          confirmInput = 3'd6;

always@(*)
begin
    case(S)
        START: 
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = START;
        end
        firstChoice:
        begin
            //if (userInput == 1'b1)
                //NS = confirmInput;
            //else    
                NS = firstChoice;
        end
        secondChoice:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = secondChoice;
        end
        thirdChoice:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = thirdChoice;
        end
        fourthChoice:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = fourthChoice;
        end
        ending:
        begin
            if (userInput == 1'b1)
                NS = confirmInput;
            else    
                NS = ending;
        end
        confirmInput:
        begin
            if (userInput == 1'b0)
            begin
                case(LS)
                    START: NS = firstChoice;
                    firstChoice: NS = secondChoice;
                    secondChoice: NS = thirdChoice;
                    thirdChoice: NS = fourthChoice;
                    fourthChoice: NS = ending;
                    ending: NS = START;
                endcase
            end
            else
                NS = confirmInput;
        end
    endcase
end

always@(posedge clk or negedge rst)
begin
    if (rst == 1'b0)
    begin
        frame <= 1344'b011000000001000001011000001000011100001100000010010001100010011000111010001100101101000011100001001000110001111000101110000000000110001111111000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110;
    end
        case(S)
            START:
            begin
                frame <= 1344'b011000000001000001011000001000011100001100000010010001100010011000111010001100101101000011100001001000110001111000101110000000000110001111111000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110;
                LS <= START;
            end
            firstChoice:
            begin
                frame <= 1344'b011001000011100010100100011000000000010001000010010001100001111000101100000000011000000100000011010000110100011000111000001110001010000011010010011000010000100010010010001001100100010001000000101000001001000110011011010001100010110000011100001000001101100001010001100010010001010000000110000011000010000011010001011001100010000101000110001100000011100010100100011000100010000100000001000001000001000001010100001001000110000000000011011000110000010000011000000000000100000010111000110000010100011100010001100011000111010010001011111010001100100011000000000011000001000000010000100100001110000110110001100000010000111000011010010011000000000010000001101000100000011010000110100011000110000001110001010000100011000110000010100010000001101000000000010111000110000010000101110000000000110001111101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110100011010001101000110;
            end
        endcase
end

always@(*)
begin
    case(choice)
    4'b1110:
    begin
        userInput = 1'b1;
        selection = 8'd1;
    end
    4'b1101:
    begin
        userInput = 1'b1;
        selection = 8'd2;
    end
    4'b1011:
    begin
        userInput = 1'b1;
        selection = 8'd3;
    end
    4'b0111:
    begin
        userInput = 1'b1;
        selection = 8'd4;
    end
    default:
    begin
        userInput = 1'b0;
        selection = 8'd0;
    end
    endcase
end

endmodule